module PC_adder (
     input [31:0] a,b,
     input[31:0] c
);
   assign c=a+b;  
endmodule